--Filename: letters_pak.vhd
--
--Description: 
--Letters package, allows the use of 'a' to 'z' in the code,
--rather than forcing binary representations
--Will also handle conversion functions into and out of the letters type
--
--
--    Copyright (C) 2013 Stephen Jeapes (vhdl-enigma@arcoarena.co.uk)
--
--    This program is free software: you can redistribute it and/or modify
--    it under the terms of the GNU General Public License as published by
--    the Free Software Foundation, either version 3 of the License, or
--    (at your option) any later version.
--
--    This program is distributed in the hope that it will be useful,
--    but WITHOUT ANY WARRANTY; without even the implied warranty of
--    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--    GNU General Public License for more details.
--
--    You should have received a copy of the GNU General Public License
--    along with this program.  If not, see <http://www.gnu.org/licenses/>.




package letters_pak is

type letter is (a,b,c,d,e,f,g,h,i,j,k,l,m,n,o,p,q,r,s,t,u,v,w,x,y,z,' '); --! An enumerated type for letters of the alphabet, purely for readability
type letter_mapping is array(letter) of letter; --! An array type used to map the incoming letter to an outgoing letter

type wheel_variants is ('1','2','3','4','5','6','7','8',beta,gamma); --! The wheel types available
type wheel_order is array(3 downto 0) of wheel_variants; --! The wheels fitted in the machine, highest wheel number to lowest, if only 3 wheels are used the MSB will be ignored

end letters_pak;

package body letters_pak is



end letters_pak;
